-- VHDL model created from schematic schema.sch -- Feb 14 10:00:37 2019

library IEEE;
use IEEE.std_logic_1164.all;
library xp2;
use xp2.components.all;

entity SCHEMA is
end SCHEMA;

architecture SCHEMATIC of SCHEMA is

   SIGNAL gnd : std_logic := '0';
   SIGNAL vcc : std_logic := '1';


begin


end SCHEMATIC;
