-- VHDL model created from schematic a.sch -- May 09 10:40:02 2019

library IEEE;
use IEEE.std_logic_1164.all;
library xp2;
use xp2.components.all;

entity A is
end A;

architecture SCHEMATIC of A is

   SIGNAL gnd : std_logic := '0';
   SIGNAL vcc : std_logic := '1';


begin


end SCHEMATIC;
